package i2c_types_pkg;

typedef enum bit {I2_WRITE=1'b0, I2_READ=1'b1} i2c_op_t;

endpackage