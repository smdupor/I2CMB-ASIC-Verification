
//asdfasdfasdfasdfasdfasdfasdfasdf  




