package i2cmb_env_pkg;

`include "src/i2cmb_coverage.svh"
`include "src/i2cmb_env_configuration.svh"
`include "src/i2cmb_generator.svh"
`include "src/i2cmb_predictor.svh"
`include "src/i2cmb_scoreboard.svh"
`include "src/i2cmb_test.svh"


endpackage